package polara_pkg;
	`include "axi/assign.svh"
    `include "axi/typedef.svh"
    `include "common_cells/registers.svh"
endpackage : polara_pkg