package polara_pkg;
	
endpackage : polara_pkg