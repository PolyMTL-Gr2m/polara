package polara_pkg;
	`include "axi/assign.svh"
    `include "axi/typedef.svh"
    `include "register_typedef.svh"
endpackage : polara_pkg